module SIPO_test;
  reg clk;
  reg reset;
  reg in;
  wire [7:0] count;
  wire frame;
  wire [3:0] out;
  wire flag;

 ini d1(clk,reset,count,frame,out,in,flag);
  initial
    begin
      in = 1'b0;
      clk = 1'b1;
      reset = 1'b1;
      #10 reset= 1'b0;

      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #5 in = 1'b0;
      #5 in = 1'b1;
      #10 in = 1'b1;
      #5 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;

      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b0;

      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b1;
      #10 in = 1'b0;
      #10 in = 1'b0;
      #10 in = 1'b1;


  
   end
   always #10 clk = ~clk;
 initial
   #100000 $finish;
 endmodule

